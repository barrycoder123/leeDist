library ieee;

package array_pkg is 
    type array_type is array(3 downto 0) of unsigned (3 downto 0);
end package array_pkg;
