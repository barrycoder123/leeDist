library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity leeDist is 

    port (



         );


end leeDist;


architecture data_flow of leeDist is 


begin 




end data_flow;
